module convolution(
    input clk,
    input rst,
    input start,
    input [6:0] X,
    input [6:0] Y,
    input [6:0] Z,
    output done);

    wire is_finished, co_row_filter, co_temp_y, co_temp_x, co_y3, co_mac, co_buf_mac_index, co_shift;
    wire load_addrs, load_row_img, init_counters, row_img_en, col_img_en, row_filter_en, row_res_en ,init_temps_counter;
    wire sel_mem_w, buf8_we, buf4w_we, buf4f_we, shift_en, y_load_buf8_e, x_load_buf8_e, mac_c_en, macbuf_c_en;
    wire shift_c_en, jump, c3_en, load_mac, init_mac, en_mac_c, step_c_en, init_mac_buf, buf_mac_we, we_memory;
    wire load_row_img_temp, row_img_temp_en;

    controller cntrl( 
        .clk(clk), 
        .rst(rst), 
        .start(start), 
        .is_finished(is_finished), 
        .co_row_filter(co_row_filter), 
        .co_temp_y(co_temp_y), 
        .co_temp_x(co_temp_x), 
        .co_y3(co_y3), 
        .co_mac(co_mac),
        .co_buf_mac_index(co_buf_mac_index), 
        .co_shift(co_shift), 
        .load_addrs(load_addrs), 
        .load_row_img(load_row_img), 
        .init_counters(init_counters),
        .init_temps_counter(init_temps_counter), 
        .row_img_en(row_img_en),
        .col_img_en(col_img_en),
        .load_row_img_temp(load_row_img_temp),
        .row_img_temp_en(row_img_temp_en), 
        .row_filter_en(row_filter_en), 
        .row_res_en(row_res_en), 
        .sel_mem_w(sel_mem_w), 
        .buf8_we(buf8_we), 
        .buf4w_we(buf4w_we), 
        .buf4f_we(buf4f_we),
        .shift_en(shift_en), 
        .y_load_buf8_e(y_load_buf8_e), 
        .x_load_buf8_e(x_load_buf8_e), 
        .mac_c_en(mac_c_en), 
        .macbuf_c_en(macbuf_c_en), 
        .shift_c_en(shift_c_en), 
        .jump(jump),
        .c3_en(c3_en), 
        .load_mac(load_mac), 
        .init_mac(init_mac), 
        .en_mac_c(en_mac_c), 
        .step_c_en(step_c_en), 
        .init_mac_buf(init_mac_buf), 
        .buf_mac_we(buf_mac_we), 
        .we_memory(we_memory), 
        .done(done)
    );

    datapath dp( 
        .clk(clk), 
        .load_addrs(load_addrs), 
        .load_row_img(load_row_img), 
        .init_counters(init_counters), 
        .init_temps_counter(init_temps_counter), 
        .row_img_en(row_img_en), 
        .col_img_en(col_img_en), 
        .load_row_img_temp(load_row_img_temp),
        .row_img_temp_en(row_img_temp_en),
        .row_filter_en(row_filter_en), 
        .row_res_en(row_res_en), 
        .sel_mem_w(sel_mem_w), 
        .buf8_we(buf8_we), 
        .buf4w_we(buf4w_we), 
        .buf4f_we(buf4f_we), 
        .buf16_she(shift_en), 
        .y_load_buf8_e(y_load_buf8_e), 
        .x_load_buf8_e(x_load_buf8_e), 
        .mac_c_en(mac_c_en), 
        .jump(jump), 
        .c3_en(c3_en), 
        .load_mac(load_mac), 
        .init_mac(init_mac), 
        .en_mac_c(en_mac_c), 
        .step_c_en(step_c_en), 
        .init_mac_buf(init_mac_buf), 
        .buf_mac_we(buf_mac_we), 
        .we_memory(we_memory), 
        .macbuf_c_en(macbuf_c_en), 
        .shift_c_en(shift_c_en), 
        .X(X), 
        .Y(Y), 
        .Z(Z), 
        .co_steps(is_finished), 
        .co_row_filter(co_row_filter), 
        .co_temp_y(co_temp_y), 
        .co_temp_x(co_temp_x), 
        .co_y3(co_y3), 
        .co_mac(co_mac), 
        .co_buf_mac_index(co_buf_mac_index), 
        .co_shift(co_shift)
    );

endmodule
