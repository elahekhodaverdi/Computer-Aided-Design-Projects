`timescale 1ps/1ps

module encoder #(parameter ) (
    ports
);
    
endmodule