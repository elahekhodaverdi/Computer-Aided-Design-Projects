module dp ();
    
endmodule