module check (a, is_finished);
    input [3:0] a;
    output is_finished;
    AND()
    
endmodule