module AND(a, b , out);
    input a, b;
    output out;
    

endmodule